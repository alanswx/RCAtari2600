library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity barnstorming is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of barnstorming is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"78",X"D8",X"A2",X"00",X"A9",X"00",X"95",X"00",X"9A",X"E8",X"D0",X"FA",X"20",X"47",X"FD",X"A5",
		X"82",X"D0",X"08",X"A2",X"01",X"86",X"82",X"CA",X"4C",X"4F",X"F6",X"A2",X"07",X"BD",X"AD",X"F0",
		X"45",X"85",X"25",X"86",X"95",X"87",X"E0",X"01",X"B0",X"02",X"95",X"09",X"CA",X"10",X"EE",X"A9",
		X"21",X"A2",X"00",X"20",X"BD",X"FD",X"A9",X"28",X"E8",X"86",X"0A",X"20",X"BD",X"FD",X"A5",X"DD",
		X"E8",X"20",X"BD",X"FD",X"A5",X"DD",X"18",X"69",X"40",X"C9",X"A0",X"90",X"02",X"E9",X"A0",X"E8",
		X"20",X"96",X"FD",X"85",X"02",X"85",X"2B",X"A2",X"03",X"B5",X"E8",X"20",X"9E",X"FD",X"85",X"F5",
		X"B5",X"E0",X"29",X"0F",X"05",X"F5",X"95",X"E0",X"95",X"E0",X"88",X"88",X"88",X"88",X"94",X"E4",
		X"CA",X"10",X"E6",X"A5",X"8B",X"85",X"09",X"AC",X"84",X"02",X"D0",X"FB",X"85",X"02",X"85",X"2A",
		X"84",X"01",X"84",X"04",X"84",X"05",X"A9",X"02",X"45",X"85",X"25",X"86",X"85",X"06",X"85",X"07",
		X"A2",X"01",X"85",X"02",X"85",X"2A",X"CA",X"10",X"F9",X"A0",X"07",X"85",X"02",X"85",X"2A",X"B1",
		X"92",X"85",X"1B",X"B1",X"94",X"85",X"1C",X"88",X"10",X"F1",X"4C",X"F1",X"F0",X"D6",X"00",X"D0",
		X"1A",X"88",X"0E",X"14",X"12",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",
		X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"D0",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"D0",X"D6",X"FF",X"FF",X"EE",X"88",X"00",X"00",X"00",X"00",X"10",X"15",X"15",
		X"25",X"85",X"02",X"85",X"2A",X"C8",X"84",X"1B",X"84",X"1C",X"C8",X"84",X"05",X"A0",X"03",X"84",
		X"04",X"EA",X"85",X"F9",X"85",X"10",X"85",X"11",X"A2",X"01",X"85",X"02",X"85",X"2A",X"A0",X"00",
		X"85",X"F9",X"C6",X"F5",X"A9",X"07",X"85",X"F5",X"A5",X"BB",X"C9",X"50",X"CA",X"85",X"2B",X"10",
		X"E9",X"90",X"05",X"84",X"04",X"84",X"05",X"CA",X"86",X"F7",X"A4",X"F5",X"B1",X"B9",X"19",X"D7",
		X"FD",X"25",X"F7",X"85",X"1B",X"B1",X"BB",X"85",X"1C",X"85",X"02",X"85",X"2A",X"B1",X"C1",X"85",
		X"F6",X"B1",X"BF",X"AA",X"B1",X"BD",X"19",X"DC",X"FD",X"A4",X"F6",X"85",X"1B",X"86",X"1C",X"84",
		X"1B",X"C6",X"F5",X"10",X"D5",X"85",X"02",X"85",X"2A",X"A9",X"00",X"85",X"1B",X"85",X"1C",X"4C",
		X"70",X"F1",X"14",X"14",X"0E",X"14",X"14",X"0E",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",
		X"A2",X"0C",X"BD",X"93",X"FF",X"45",X"85",X"25",X"86",X"E0",X"08",X"B0",X"1C",X"85",X"02",X"85",
		X"2A",X"85",X"09",X"A5",X"8E",X"85",X"08",X"BD",X"E5",X"F0",X"85",X"0D",X"BD",X"E4",X"FD",X"85",
		X"0E",X"BD",X"EC",X"FD",X"85",X"0F",X"4C",X"9F",X"F1",X"85",X"02",X"85",X"2A",X"85",X"09",X"CA",
		X"10",X"D0",X"A2",X"00",X"A4",X"87",X"A5",X"8A",X"85",X"02",X"85",X"2A",X"85",X"08",X"84",X"09",
		X"86",X"0D",X"86",X"0E",X"86",X"0F",X"86",X"05",X"86",X"0A",X"A5",X"89",X"85",X"11",X"85",X"07",
		X"A9",X"F0",X"85",X"21",X"85",X"02",X"85",X"2A",X"20",X"BC",X"FD",X"20",X"BC",X"FD",X"85",X"2B",
		X"A2",X"04",X"86",X"DB",X"A4",X"8F",X"85",X"02",X"85",X"2A",X"C0",X"15",X"B0",X"29",X"B1",X"9A",
		X"85",X"1C",X"B9",X"45",X"FF",X"85",X"0E",X"CA",X"86",X"DB",X"B5",X"E0",X"85",X"04",X"85",X"EC",
		X"A9",X"00",X"85",X"0E",X"88",X"C0",X"15",X"B0",X"19",X"B1",X"9A",X"85",X"1C",X"B9",X"45",X"FF",
		X"84",X"F5",X"85",X"0E",X"4C",X"1B",X"F2",X"A9",X"00",X"85",X"0E",X"85",X"1C",X"85",X"F9",X"4C",
		X"E7",X"F1",X"A9",X"00",X"85",X"0E",X"85",X"1C",X"4C",X"00",X"F2",X"85",X"02",X"85",X"2A",X"B5",
		X"E4",X"AA",X"30",X"21",X"E0",X"05",X"B0",X"49",X"E0",X"02",X"B0",X"29",X"CA",X"10",X"FD",X"EA",
		X"85",X"10",X"20",X"BC",X"FD",X"A9",X"00",X"85",X"0E",X"88",X"C0",X"15",X"B0",X"04",X"B1",X"9A",
		X"85",X"1C",X"4C",X"91",X"F2",X"85",X"F9",X"85",X"F9",X"85",X"F9",X"8D",X"10",X"00",X"A9",X"60",
		X"85",X"20",X"4C",X"32",X"F2",X"85",X"F9",X"CA",X"CA",X"85",X"F9",X"CA",X"10",X"FD",X"8D",X"10",
		X"00",X"A9",X"00",X"85",X"0E",X"88",X"C0",X"15",X"B0",X"04",X"B1",X"9A",X"85",X"1C",X"4C",X"91",
		X"F2",X"E9",X"05",X"AA",X"88",X"C0",X"15",X"90",X"07",X"85",X"F9",X"C6",X"F5",X"4C",X"85",X"F2",
		X"B1",X"9A",X"EA",X"85",X"1C",X"A9",X"00",X"85",X"0E",X"85",X"F9",X"CA",X"10",X"FD",X"8D",X"10",
		X"00",X"85",X"02",X"85",X"2A",X"C0",X"15",X"90",X"06",X"EA",X"85",X"F9",X"4C",X"A4",X"F2",X"B9",
		X"45",X"FF",X"85",X"0E",X"A6",X"DB",X"F0",X"60",X"AD",X"F1",X"00",X"85",X"9C",X"A5",X"EC",X"85",
		X"20",X"A5",X"8C",X"8D",X"06",X"00",X"A2",X"0C",X"A5",X"DE",X"85",X"0E",X"88",X"C0",X"15",X"B0",
		X"3A",X"B1",X"9A",X"85",X"1C",X"B9",X"45",X"FF",X"85",X"0E",X"84",X"F5",X"8A",X"A8",X"85",X"2A",
		X"A6",X"DB",X"B5",X"ED",X"85",X"9C",X"B1",X"9C",X"85",X"1B",X"98",X"AA",X"A4",X"F5",X"A5",X"07",
		X"85",X"F9",X"85",X"2B",X"CA",X"10",X"D1",X"A2",X"00",X"86",X"EC",X"86",X"0E",X"A6",X"DB",X"88",
		X"05",X"02",X"15",X"B1",X"95",X"B1",X"85",X"2C",X"4C",X"D6",X"F1",X"85",X"1C",X"84",X"F5",X"8A",
		X"A8",X"EA",X"EA",X"EA",X"EA",X"4C",X"CE",X"F2",X"A5",X"EC",X"85",X"20",X"85",X"F9",X"85",X"F9",
		X"A2",X"47",X"88",X"C0",X"15",X"B0",X"13",X"A9",X"00",X"85",X"0E",X"B1",X"9A",X"85",X"1C",X"B9",
		X"45",X"FF",X"EA",X"EA",X"EA",X"85",X"0E",X"4C",X"30",X"F3",X"A9",X"00",X"85",X"0E",X"85",X"1C",
		X"85",X"02",X"85",X"2A",X"20",X"BA",X"FD",X"20",X"BC",X"FD",X"85",X"2B",X"A9",X"00",X"85",X"0E",
		X"E6",X"F5",X"C6",X"F5",X"88",X"C0",X"15",X"B0",X"0C",X"B1",X"9A",X"85",X"1C",X"B9",X"45",X"FF",
		X"85",X"0E",X"4C",X"5E",X"F3",X"A9",X"00",X"85",X"1C",X"85",X"0E",X"4C",X"5E",X"F3",X"85",X"02",
		X"85",X"2A",X"A5",X"F3",X"D0",X"46",X"20",X"BC",X"FD",X"A5",X"89",X"85",X"06",X"EA",X"EA",X"EA",
		X"EA",X"88",X"A9",X"00",X"85",X"0E",X"C0",X"15",X"90",X"07",X"84",X"F5",X"8A",X"A8",X"4C",X"90",
		X"F3",X"B1",X"9A",X"85",X"1C",X"B9",X"45",X"FF",X"84",X"F5",X"86",X"F6",X"A4",X"F6",X"85",X"0E",
		X"85",X"02",X"85",X"2A",X"E0",X"39",X"B0",X"06",X"B9",X"5A",X"FF",X"4C",X"A0",X"F3",X"B1",X"A6",
		X"25",X"F4",X"85",X"1B",X"A4",X"F5",X"CA",X"10",X"C8",X"4C",X"83",X"F4",X"20",X"B9",X"FD",X"EA",
		X"EA",X"85",X"F9",X"88",X"A9",X"00",X"85",X"0E",X"C0",X"15",X"90",X"09",X"85",X"1C",X"84",X"F5",
		X"8A",X"A8",X"4C",X"D4",X"F3",X"B1",X"9A",X"85",X"1C",X"B9",X"45",X"FF",X"84",X"F5",X"86",X"F6",
		X"A4",X"F6",X"85",X"0E",X"85",X"02",X"85",X"2A",X"A5",X"8C",X"85",X"06",X"B9",X"01",X"FF",X"25",
		X"F4",X"85",X"1B",X"A4",X"F5",X"EA",X"EA",X"EA",X"E0",X"30",X"F0",X"1E",X"CA",X"10",X"C4",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"85",X"1C",X"84",X"F5",X"4C",X"20",X"F4",X"CA",X"88",X"A9",X"00",X"85",X"0E",
		X"C0",X"15",X"B0",X"EF",X"B1",X"9A",X"85",X"1C",X"B9",X"45",X"FF",X"84",X"F5",X"EA",X"85",X"0E",
		X"8A",X"A8",X"A9",X"07",X"85",X"02",X"85",X"2A",X"85",X"04",X"B9",X"B5",X"F0",X"45",X"85",X"25",
		X"86",X"85",X"06",X"A5",X"A2",X"85",X"1B",X"A4",X"F5",X"CA",X"E0",X"18",X"B0",X"CD",X"A9",X"E0",
		X"85",X"20",X"88",X"A9",X"00",X"85",X"0E",X"C0",X"15",X"B0",X"2D",X"B1",X"9A",X"85",X"1C",X"B9",
		X"45",X"FF",X"84",X"F5",X"85",X"0E",X"8A",X"A8",X"A9",X"07",X"EA",X"85",X"2A",X"85",X"04",X"B9",
		X"B5",X"F0",X"45",X"85",X"25",X"86",X"85",X"06",X"A5",X"A3",X"85",X"1B",X"A4",X"F5",X"85",X"2B",
		X"85",X"F9",X"CA",X"10",X"CD",X"4C",X"83",X"F4",X"85",X"1C",X"84",X"F5",X"EA",X"EA",X"EA",X"EA",
		X"4C",X"56",X"F4",X"A5",X"07",X"05",X"02",X"05",X"B1",X"85",X"B1",X"85",X"2C",X"85",X"02",X"85",
		X"2A",X"A9",X"00",X"85",X"1C",X"85",X"1B",X"A5",X"89",X"85",X"09",X"A5",X"8C",X"85",X"06",X"85",
		X"07",X"A9",X"06",X"85",X"04",X"85",X"05",X"A0",X"0C",X"C0",X"07",X"A2",X"00",X"B0",X"02",X"A2",
		X"02",X"85",X"02",X"85",X"2A",X"86",X"1D",X"86",X"1E",X"B9",X"62",X"F1",X"45",X"85",X"25",X"86",
		X"85",X"09",X"88",X"10",X"E4",X"A0",X"02",X"A9",X"00",X"A6",X"8D",X"85",X"02",X"85",X"2A",X"85",
		X"1D",X"85",X"1E",X"86",X"09",X"88",X"10",X"EF",X"85",X"02",X"85",X"2A",X"A5",X"88",X"85",X"09",
		X"85",X"02",X"85",X"2A",X"85",X"F9",X"A2",X"00",X"86",X"2B",X"86",X"0B",X"86",X"0C",X"E8",X"86",
		X"04",X"85",X"F9",X"85",X"10",X"85",X"11",X"E8",X"E8",X"86",X"05",X"A9",X"10",X"85",X"21",X"A0",
		X"07",X"B1",X"96",X"85",X"F5",X"85",X"02",X"85",X"2A",X"B9",X"58",X"FE",X"85",X"1B",X"B9",X"60",
		X"FE",X"85",X"1C",X"EA",X"B9",X"70",X"FE",X"AA",X"B9",X"68",X"FE",X"85",X"1B",X"86",X"1C",X"A5",
		X"F5",X"85",X"1C",X"85",X"2B",X"88",X"10",X"D9",X"C8",X"84",X"1B",X"84",X"1C",X"A9",X"21",X"A2",
		X"82",X"85",X"02",X"8D",X"96",X"02",X"86",X"01",X"A9",X"FE",X"85",X"93",X"85",X"95",X"85",X"97",
		X"A5",X"D3",X"29",X"F0",X"4A",X"D0",X"02",X"A9",X"50",X"85",X"92",X"A6",X"80",X"E8",X"8A",X"0A",
		X"0A",X"0A",X"85",X"96",X"A5",X"D3",X"29",X"0F",X"0A",X"0A",X"0A",X"85",X"94",X"A0",X"08",X"A2",
		X"02",X"B5",X"B5",X"29",X"0F",X"0A",X"0A",X"0A",X"99",X"B9",X"00",X"CA",X"30",X"0E",X"88",X"88",
		X"B5",X"B6",X"29",X"F0",X"4A",X"99",X"B9",X"00",X"88",X"88",X"10",X"E5",X"D8",X"A5",X"D1",X"D0",
		X"04",X"A5",X"A8",X"30",X"00",X"A5",X"81",X"29",X"07",X"D0",X"0E",X"A6",X"DC",X"E8",X"8A",X"29",
		X"07",X"85",X"DC",X"A8",X"B9",X"BA",X"FE",X"85",X"F1",X"A0",X"00",X"A5",X"81",X"29",X"01",X"D0",
		X"02",X"A0",X"20",X"84",X"F2",X"A2",X"05",X"A0",X"00",X"A5",X"A8",X"C9",X"20",X"B0",X"06",X"A5",
		X"D1",X"D0",X"02",X"B4",X"C9",X"94",X"15",X"CA",X"10",X"ED",X"A5",X"AB",X"D0",X"0E",X"A5",X"D6",
		X"C9",X"0A",X"B0",X"08",X"A5",X"8F",X"C9",X"7D",X"B0",X"02",X"E6",X"8F",X"AD",X"84",X"02",X"D0",
		X"FB",X"A0",X"82",X"84",X"02",X"84",X"00",X"84",X"02",X"84",X"02",X"84",X"02",X"85",X"00",X"E6",
		X"81",X"D0",X"07",X"E6",X"A8",X"D0",X"03",X"38",X"66",X"A8",X"A0",X"FF",X"AD",X"82",X"02",X"29",
		X"08",X"D0",X"02",X"A0",X"0F",X"98",X"A0",X"00",X"24",X"A8",X"10",X"04",X"29",X"F7",X"A4",X"A8",
		X"84",X"85",X"06",X"85",X"85",X"86",X"A9",X"30",X"85",X"02",X"8D",X"96",X"02",X"AD",X"80",X"02",
		X"A8",X"A6",X"AC",X"F0",X"02",X"A0",X"0F",X"98",X"4A",X"4A",X"4A",X"4A",X"85",X"84",X"C8",X"F0",
		X"07",X"A9",X"00",X"85",X"A8",X"4C",X"2C",X"F6",X"24",X"0C",X"10",X"F5",X"AD",X"82",X"02",X"4A",
		X"B0",X"05",X"A2",X"A8",X"4C",X"04",X"F0",X"A0",X"00",X"4A",X"B0",X"2F",X"A5",X"83",X"F0",X"04",
		X"C6",X"83",X"10",X"29",X"E6",X"80",X"A5",X"80",X"C9",X"03",X"D0",X"03",X"20",X"CA",X"FD",X"A5",
		X"80",X"29",X"03",X"85",X"80",X"85",X"A8",X"A9",X"AA",X"85",X"D3",X"85",X"B5",X"85",X"B6",X"85",
		X"B7",X"85",X"B8",X"A9",X"50",X"85",X"BB",X"A0",X"1E",X"84",X"D1",X"84",X"83",X"A5",X"A8",X"30",
		X"04",X"A5",X"D1",X"F0",X"03",X"4C",X"1B",X"F0",X"A5",X"CF",X"D0",X"0D",X"24",X"0C",X"10",X"03",
		X"4C",X"1B",X"F0",X"A9",X"01",X"85",X"CF",X"85",X"81",X"24",X"B0",X"10",X"3C",X"A5",X"EB",X"05",
		X"E9",X"05",X"EA",X"D0",X"0C",X"A5",X"8F",X"C9",X"7D",X"D0",X"06",X"A9",X"C2",X"85",X"9A",X"E6",
		X"D1",X"A5",X"81",X"A6",X"D6",X"F0",X"13",X"E0",X"1A",X"B0",X"09",X"29",X"03",X"D0",X"0B",X"C6",
		X"D6",X"4C",X"BA",X"F6",X"29",X"01",X"D0",X"02",X"C6",X"D6",X"A5",X"81",X"29",X"03",X"D0",X"06",
		X"A5",X"D4",X"F0",X"02",X"C6",X"D4",X"4C",X"56",X"F7",X"A5",X"B5",X"C9",X"05",X"D0",X"05",X"E6",
		X"D1",X"4C",X"56",X"F7",X"18",X"A5",X"B8",X"69",X"AB",X"85",X"B8",X"A9",X"01",X"F8",X"65",X"B7",
		X"85",X"B7",X"A5",X"B6",X"69",X"00",X"85",X"B6",X"D8",X"C9",X"60",X"90",X"06",X"A9",X"00",X"85",
		X"B6",X"E6",X"B5",X"A5",X"81",X"29",X"01",X"D0",X"31",X"24",X"0C",X"30",X"16",X"A6",X"D6",X"E8",
		X"E0",X"25",X"90",X"02",X"A2",X"25",X"86",X"D6",X"A5",X"81",X"29",X"07",X"D0",X"02",X"E6",X"D4",
		X"4C",X"2A",X"F7",X"A5",X"81",X"29",X"07",X"D0",X"02",X"C6",X"D4",X"A6",X"D6",X"E0",X"18",X"B0",
		X"05",X"E6",X"D6",X"4C",X"2A",X"F7",X"F0",X"02",X"C6",X"D6",X"A5",X"D4",X"10",X"02",X"A9",X"00",
		X"C9",X"08",X"90",X"02",X"A9",X"07",X"85",X"D4",X"A2",X"00",X"A5",X"81",X"29",X"01",X"D0",X"16",
		X"A5",X"84",X"49",X"0F",X"29",X"03",X"F0",X"0C",X"A5",X"D5",X"18",X"69",X"05",X"C9",X"17",X"90",
		X"02",X"A9",X"17",X"AA",X"86",X"D5",X"EA",X"A5",X"D0",X"A2",X"03",X"85",X"F5",X"29",X"01",X"F0",
		X"7D",X"B5",X"E8",X"D0",X"02",X"A9",X"A0",X"A4",X"D8",X"88",X"84",X"F6",X"38",X"E5",X"F6",X"85",
		X"F7",X"F0",X"29",X"C9",X"A1",X"B0",X"25",X"B5",X"E0",X"29",X"F0",X"95",X"E0",X"B4",X"C5",X"A5",
		X"F7",X"D9",X"06",X"FD",X"B0",X"56",X"B5",X"E0",X"15",X"C5",X"95",X"E0",X"A5",X"F7",X"4C",X"DC",
		X"F7",X"B5",X"E0",X"15",X"C5",X"95",X"E0",X"A5",X"F7",X"4C",X"DC",X"F7",X"B5",X"E0",X"29",X"0F",
		X"C9",X"00",X"F0",X"13",X"A8",X"B9",X"01",X"FD",X"95",X"E8",X"B5",X"E0",X"29",X"F0",X"95",X"E0",
		X"A9",X"00",X"95",X"C5",X"4C",X"DE",X"F7",X"F6",X"C2",X"B5",X"C2",X"29",X"03",X"95",X"C2",X"A8",
		X"86",X"F8",X"A6",X"80",X"A9",X"FD",X"85",X"99",X"BD",X"EC",X"FC",X"85",X"98",X"B1",X"98",X"A6",
		X"F8",X"95",X"C5",X"BD",X"F0",X"FC",X"45",X"D0",X"85",X"D0",X"A9",X"00",X"95",X"E8",X"A5",X"F5",
		X"4A",X"CA",X"F0",X"03",X"4C",X"5B",X"F7",X"A5",X"D1",X"D0",X"3C",X"A5",X"81",X"29",X"01",X"D0",
		X"0C",X"24",X"0C",X"10",X"06",X"A5",X"81",X"29",X"03",X"D0",X"02",X"E6",X"90",X"A6",X"90",X"E0",
		X"03",X"90",X"04",X"A2",X"00",X"86",X"90",X"BD",X"78",X"FE",X"85",X"9A",X"A5",X"81",X"29",X"03",
		X"D0",X"02",X"E6",X"91",X"A6",X"91",X"E0",X"03",X"90",X"02",X"A2",X"00",X"86",X"91",X"BD",X"D7",
		X"FE",X"85",X"A6",X"A9",X"FF",X"85",X"A7",X"A6",X"AB",X"F0",X"03",X"CA",X"86",X"AB",X"A6",X"D2",
		X"F0",X"03",X"CA",X"86",X"D2",X"A2",X"03",X"A5",X"F1",X"95",X"ED",X"CA",X"D0",X"F9",X"86",X"CE",
		X"A9",X"1F",X"38",X"E5",X"D4",X"85",X"CB",X"A9",X"0A",X"85",X"C9",X"A5",X"81",X"29",X"03",X"D0",
		X"0C",X"E6",X"A9",X"A5",X"A9",X"C9",X"03",X"90",X"02",X"A9",X"03",X"85",X"A9",X"A5",X"A9",X"A8",
		X"24",X"0C",X"30",X"01",X"C8",X"84",X"CD",X"A4",X"A4",X"A9",X"FC",X"85",X"99",X"A6",X"80",X"BD",
		X"E4",X"FC",X"85",X"98",X"B1",X"98",X"85",X"F5",X"A5",X"E8",X"C9",X"40",X"B0",X"1D",X"A0",X"0A",
		X"84",X"CA",X"A0",X"15",X"84",X"CC",X"C9",X"20",X"90",X"04",X"C6",X"CC",X"49",X"3F",X"4A",X"A4",
		X"8F",X"C0",X"55",X"90",X"02",X"A9",X"00",X"25",X"F4",X"85",X"CE",X"A6",X"AC",X"F0",X"06",X"CA",
		X"86",X"AC",X"4C",X"03",X"F9",X"CA",X"86",X"AA",X"24",X"B1",X"30",X"03",X"4C",X"99",X"F9",X"A5",
		X"F5",X"4A",X"B0",X"48",X"A5",X"DF",X"38",X"E9",X"18",X"C9",X"22",X"B0",X"08",X"A9",X"01",X"85",
		X"CD",X"A9",X"00",X"85",X"CE",X"A5",X"DF",X"C9",X"0C",X"90",X"11",X"A9",X"64",X"2C",X"82",X"02",
		X"50",X"02",X"A9",X"79",X"85",X"F8",X"A5",X"8F",X"C5",X"F8",X"90",X"20",X"A4",X"D2",X"D0",X"18",
		X"A9",X"50",X"85",X"D2",X"A5",X"DF",X"C9",X"30",X"90",X"0E",X"A5",X"D3",X"F0",X"0A",X"F8",X"38",
		X"E9",X"01",X"85",X"D3",X"D0",X"02",X"C6",X"B0",X"D8",X"4C",X"99",X"F9",X"A9",X"46",X"85",X"AB",
		X"4A",X"85",X"AC",X"A9",X"08",X"85",X"CA",X"A2",X"00",X"86",X"CD",X"86",X"D4",X"86",X"B1",X"A5",
		X"AC",X"4A",X"85",X"CE",X"A5",X"AA",X"30",X"3E",X"A5",X"8F",X"A6",X"AA",X"E0",X"01",X"F0",X"12",
		X"18",X"69",X"04",X"AA",X"A5",X"81",X"29",X"01",X"D0",X"05",X"8A",X"38",X"E9",X"09",X"AA",X"4C",
		X"48",X"F9",X"18",X"69",X"05",X"AA",X"A5",X"81",X"29",X"01",X"D0",X"0C",X"8A",X"38",X"E9",X"06",
		X"C9",X"64",X"B0",X"03",X"18",X"69",X"02",X"AA",X"86",X"8F",X"A5",X"AA",X"30",X"08",X"F0",X"26",
		X"4A",X"B0",X"14",X"4C",X"8B",X"F9",X"A5",X"F5",X"4A",X"B0",X"2A",X"A5",X"DF",X"C9",X"39",X"B0",
		X"2A",X"A5",X"8F",X"C9",X"5A",X"90",X"0F",X"A9",X"01",X"85",X"AA",X"A9",X"01",X"85",X"D8",X"A9",
		X"04",X"85",X"D6",X"4C",X"99",X"F9",X"A9",X"01",X"85",X"D8",X"A9",X"04",X"85",X"D6",X"A9",X"00",
		X"85",X"AA",X"4C",X"99",X"F9",X"A5",X"E8",X"C9",X"20",X"90",X"EB",X"A2",X"00",X"86",X"D6",X"CA",
		X"86",X"D8",X"A9",X"02",X"85",X"AA",X"4C",X"99",X"F9",X"A2",X"03",X"B4",X"AC",X"F0",X"26",X"88",
		X"94",X"AC",X"C0",X"27",X"90",X"0C",X"A9",X"0C",X"85",X"CA",X"A9",X"1F",X"85",X"CC",X"A9",X"05",
		X"85",X"CE",X"B4",X"E8",X"F0",X"1F",X"C8",X"C8",X"94",X"E8",X"A5",X"F2",X"95",X"ED",X"A9",X"00",
		X"95",X"B1",X"4C",X"D5",X"F9",X"B5",X"B1",X"10",X"0C",X"A9",X"00",X"85",X"D4",X"A9",X"10",X"85",
		X"D6",X"A9",X"30",X"95",X"AC",X"CA",X"D0",X"C3",X"A2",X"01",X"A5",X"AC",X"F0",X"02",X"A2",X"00",
		X"B5",X"D5",X"E0",X"01",X"D0",X"15",X"A5",X"84",X"29",X"03",X"C9",X"03",X"A5",X"D6",X"B0",X"0B",
		X"4A",X"4A",X"4A",X"4A",X"85",X"F5",X"38",X"A5",X"D6",X"E5",X"F5",X"85",X"F6",X"4A",X"4A",X"4A",
		X"4A",X"95",X"D7",X"A5",X"F6",X"29",X"0F",X"18",X"75",X"D9",X"C9",X"10",X"90",X"02",X"F6",X"D7",
		X"29",X"0F",X"95",X"D9",X"CA",X"10",X"C9",X"24",X"B0",X"30",X"2A",X"A5",X"84",X"29",X"02",X"D0",
		X"07",X"A5",X"8F",X"18",X"65",X"D7",X"85",X"8F",X"A5",X"84",X"29",X"01",X"D0",X"07",X"A5",X"8F",
		X"38",X"E5",X"D7",X"85",X"8F",X"A5",X"8F",X"C9",X"14",X"B0",X"02",X"A9",X"14",X"C9",X"7E",X"90",
		X"02",X"A9",X"7D",X"85",X"8F",X"A5",X"DD",X"38",X"E5",X"D8",X"85",X"F5",X"C9",X"A0",X"D0",X"05",
		X"A9",X"00",X"4C",X"65",X"FA",X"C9",X"F0",X"90",X"0C",X"38",X"A9",X"00",X"E5",X"F5",X"85",X"F5",
		X"38",X"A9",X"A0",X"E5",X"F5",X"85",X"DD",X"A5",X"F3",X"F0",X"17",X"38",X"A5",X"DF",X"E5",X"D8",
		X"C9",X"F0",X"90",X"04",X"A9",X"00",X"85",X"E8",X"85",X"DF",X"D0",X"03",X"4C",X"94",X"FA",X"4C",
		X"DD",X"FA",X"38",X"A5",X"E8",X"E5",X"D8",X"C9",X"F0",X"90",X"02",X"A9",X"00",X"85",X"E8",X"F0",
		X"03",X"4C",X"22",X"FB",X"A2",X"00",X"86",X"B1",X"CA",X"86",X"F4",X"E6",X"A4",X"A5",X"A4",X"29",
		X"3F",X"85",X"A4",X"A8",X"A9",X"FC",X"85",X"99",X"A6",X"80",X"BD",X"E4",X"FC",X"85",X"98",X"B1",
		X"98",X"F0",X"06",X"4A",X"B0",X"10",X"4C",X"D4",X"FA",X"A9",X"00",X"85",X"F3",X"85",X"F4",X"A9",
		X"9F",X"85",X"E8",X"4C",X"22",X"FB",X"A2",X"00",X"86",X"F3",X"CA",X"86",X"F4",X"A9",X"9F",X"85",
		X"E8",X"4C",X"22",X"FB",X"85",X"F3",X"A9",X"B7",X"85",X"DF",X"4C",X"DD",X"FA",X"A9",X"FF",X"85",
		X"A2",X"A9",X"FE",X"85",X"A3",X"A5",X"DF",X"C9",X"A0",X"90",X"08",X"E9",X"A0",X"4A",X"4A",X"AA",
		X"4C",X"06",X"FB",X"C9",X"18",X"90",X"05",X"A2",X"06",X"4C",X"06",X"FB",X"A2",X"00",X"86",X"F4",
		X"4A",X"4A",X"18",X"69",X"07",X"AA",X"A0",X"01",X"B9",X"A2",X"00",X"3D",X"F4",X"FC",X"99",X"A2",
		X"00",X"88",X"10",X"F4",X"A5",X"DF",X"38",X"E9",X"18",X"C9",X"E0",X"90",X"03",X"38",X"E9",X"60",
		X"85",X"E8",X"A6",X"D6",X"E0",X"20",X"90",X"2A",X"A9",X"3F",X"2C",X"82",X"02",X"10",X"01",X"4A",
		X"85",X"F5",X"A5",X"81",X"25",X"F5",X"D0",X"02",X"E6",X"A5",X"A5",X"A5",X"29",X"0F",X"85",X"A5",
		X"A8",X"A6",X"80",X"A9",X"FD",X"85",X"99",X"BD",X"E8",X"FC",X"85",X"98",X"B1",X"98",X"05",X"D0",
		X"85",X"D0",X"4C",X"1B",X"F0",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"03",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"00",X"03",X"02",X"03",X"03",X"03",X"02",X"03",
		X"02",X"03",X"03",X"02",X"02",X"03",X"02",X"03",X"03",X"03",X"02",X"00",X"02",X"02",X"02",X"00",
		X"02",X"02",X"02",X"00",X"02",X"02",X"03",X"00",X"03",X"03",X"03",X"02",X"02",X"02",X"03",X"02",
		X"03",X"02",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"03",
		X"03",X"03",X"02",X"02",X"03",X"03",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"02",X"02",X"03",
		X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"02",X"03",
		X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"02",X"02",X"03",
		X"03",X"02",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"03",X"02",
		X"02",X"03",X"02",X"00",X"03",X"03",X"02",X"02",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",
		X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",
		X"03",X"03",X"02",X"03",X"03",X"03",X"02",X"03",X"02",X"02",X"02",X"02",X"00",X"03",X"02",X"03",
		X"02",X"03",X"03",X"03",X"00",X"02",X"03",X"03",X"02",X"03",X"02",X"02",X"03",X"03",X"03",X"03",
		X"02",X"03",X"02",X"02",X"03",X"03",X"02",X"03",X"02",X"02",X"03",X"03",X"02",X"03",X"02",X"03",
		X"02",X"02",X"02",X"03",X"00",X"03",X"03",X"03",X"02",X"03",X"02",X"02",X"00",X"02",X"02",X"03",
		X"03",X"03",X"03",X"02",X"00",X"26",X"6C",X"AC",X"17",X"17",X"27",X"37",X"0B",X"0B",X"0F",X"13",
		X"00",X"04",X"02",X"01",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"FF",X"03",X"07",X"0F",X"1F",X"3F",
		X"7F",X"00",X"10",X"20",X"20",X"40",X"00",X"90",X"80",X"80",X"60",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"00",X"02",X"04",X"00",X"01",X"02",X"04",X"05",X"02",X"01",X"02",X"01",
		X"04",X"02",X"01",X"04",X"02",X"01",X"02",X"00",X"02",X"02",X"04",X"04",X"02",X"02",X"02",X"02",
		X"04",X"01",X"01",X"04",X"02",X"01",X"02",X"00",X"01",X"02",X"04",X"05",X"02",X"01",X"02",X"01",
		X"04",X"02",X"01",X"04",X"02",X"01",X"02",X"A9",X"00",X"85",X"9C",X"85",X"F1",X"A9",X"FF",X"85",
		X"9D",X"A9",X"C2",X"85",X"9A",X"A9",X"FE",X"85",X"9B",X"A9",X"FE",X"85",X"BA",X"85",X"BC",X"85",
		X"BE",X"85",X"C0",X"85",X"C2",X"85",X"93",X"85",X"95",X"A9",X"00",X"A6",X"80",X"E0",X"03",X"D0",
		X"04",X"A5",X"82",X"29",X"3F",X"85",X"A4",X"29",X"0F",X"85",X"A5",X"BD",X"ED",X"F0",X"85",X"D3",
		X"A9",X"7D",X"85",X"8F",X"A9",X"01",X"85",X"C3",X"85",X"C4",X"85",X"C5",X"A2",X"03",X"A9",X"00",
		X"95",X"F1",X"CA",X"10",X"F9",X"60",X"20",X"BD",X"FD",X"85",X"02",X"85",X"2A",X"60",X"18",X"69",
		X"2E",X"A8",X"29",X"0F",X"85",X"F5",X"98",X"4A",X"4A",X"4A",X"4A",X"A8",X"18",X"65",X"F5",X"C9",
		X"0F",X"90",X"03",X"E9",X"0F",X"C8",X"49",X"07",X"0A",X"0A",X"0A",X"0A",X"60",X"20",X"9E",X"FD",
		X"95",X"20",X"85",X"02",X"88",X"10",X"FD",X"95",X"10",X"60",X"A5",X"82",X"0A",X"0A",X"0A",X"45",
		X"82",X"0A",X"26",X"82",X"A5",X"82",X"60",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"0E",X"04",X"7F",X"7F",X"3F",X"0F",
		X"03",X"00",X"00",X"00",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"78",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"78",X"78",X"30",X"30",X"30",X"30",X"30",X"70",X"30",
		X"FC",X"C0",X"C0",X"78",X"0C",X"0C",X"8C",X"78",X"78",X"8C",X"0C",X"18",X"18",X"0C",X"8C",X"78",
		X"18",X"18",X"18",X"FC",X"98",X"58",X"38",X"18",X"F8",X"8C",X"0C",X"0C",X"F8",X"C0",X"C0",X"FC",
		X"78",X"CC",X"CC",X"CC",X"F8",X"C0",X"C4",X"78",X"30",X"30",X"30",X"30",X"18",X"0C",X"84",X"FC",
		X"78",X"CC",X"CC",X"78",X"78",X"CC",X"CC",X"78",X"78",X"8C",X"0C",X"7C",X"CC",X"CC",X"CC",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AD",X"A9",X"E9",X"A9",X"ED",X"41",X"0F",
		X"00",X"50",X"58",X"5C",X"56",X"53",X"11",X"F0",X"00",X"BA",X"8A",X"BA",X"A2",X"3A",X"80",X"FE",
		X"00",X"E9",X"AB",X"AF",X"AD",X"E9",X"00",X"00",X"7B",X"90",X"A5",X"00",X"04",X"0A",X"0A",X"0C",
		X"18",X"30",X"FC",X"FD",X"A1",X"40",X"11",X"21",X"08",X"31",X"65",X"B0",X"31",X"04",X"7E",X"7E",
		X"00",X"04",X"0A",X"0A",X"0C",X"18",X"30",X"FD",X"FD",X"A0",X"41",X"11",X"20",X"09",X"B1",X"64",
		X"31",X"31",X"04",X"7E",X"7E",X"00",X"04",X"0A",X"0A",X"0C",X"18",X"30",X"FD",X"FC",X"A1",X"41",
		X"10",X"21",X"09",X"30",X"E5",X"31",X"30",X"04",X"7E",X"7E",X"10",X"10",X"10",X"00",X"20",X"20",
		X"00",X"10",X"00",X"04",X"0A",X"0A",X"0C",X"18",X"30",X"FC",X"FD",X"A1",X"41",X"11",X"20",X"09",
		X"31",X"E5",X"31",X"30",X"04",X"7E",X"7E",X"6B",X"7B",X"8B",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"00",X"00",X"00",X"40",X"30",X"78",X"FC",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"78",X"FC",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"30",X"78",X"FC",X"36",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"11",X"53",X"FE",X"53",X"11",X"10",X"38",X"3C",X"3E",X"62",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"A8",X"80",X"80",X"80",X"00",X"00",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"FE",X"82",X"C6",X"82",X"AA",X"82",X"92",X"82",X"AA",X"82",X"C6",X"82",X"FE",
		X"44",X"44",X"44",X"6C",X"44",X"54",X"44",X"54",X"54",X"54",X"44",X"54",X"44",X"6C",X"44",X"44",
		X"44",X"44",X"44",X"7C",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"38",X"28",X"28",X"28",X"28",
		X"28",X"28",X"FE",X"10",X"1A",X"18",X"28",X"28",X"38",X"38",X"48",X"48",X"58",X"68",X"68",X"78",
		X"78",X"88",X"88",X"FE",X"10",X"10",X"90",X"91",X"12",X"97",X"8E",X"7F",X"8E",X"87",X"02",X"81",
		X"80",X"00",X"00",X"FE",X"10",X"10",X"90",X"11",X"92",X"97",X"0E",X"FF",X"8E",X"07",X"82",X"81",
		X"00",X"00",X"00",X"FE",X"10",X"10",X"10",X"91",X"92",X"17",X"8E",X"FF",X"0E",X"87",X"82",X"01",
		X"80",X"00",X"00",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"00",X"F0",X"00",X"F0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
